`timescale 1ns/1ns

module sim_nn_rgb;

  // define constants for multiple images
  localparam string stimuli_filenames[]  = {"training-3.ppm"};
  localparam string response_filenames[] = {"sim-training-3.ppm", "sim-training-2.ppm", "sim-gril.ppm"};
  localparam int num_files = 1;
  localparam int x_blank = 100;   // horizontal blanking
  localparam int trail = 1000;  // clock cycles after active image

  // signals of testbench
  logic clk = 0;
  logic reset_n;
  logic [2:0] enable_in;
  logic vs_in;
  logic hs_in;
  logic de_in;
  logic [7:0] r_in;
  logic [7:0] g_in;
  logic [7:0] b_in;
  logic vs_out;
  logic hs_out;
  logic de_out;
  logic [7:0] r_out;
  logic [7:0] g_out;
  logic [7:0] b_out;
  logic clk_o;
  logic [2:0] led;
  int x_size, y_size;
  int end_tb = 0;
  int mismatch = 0;

  // Clock generation
  always #20 clk = ~clk;

  // Instantiate the design under verification (DUV)
  nn_rgb duv (
    .clk(clk),
    .reset_n(reset_n),
    .enable_in(enable_in),
    .vs_in(vs_in),
    .hs_in(hs_in),
    .de_in(de_in),
    .r_in(r_in),
    .g_in(g_in),
    .b_in(b_in),
    .vs_out(vs_out),
    .hs_out(hs_out),
    .de_out(de_out),
    .r_out(r_out),
    .g_out(g_out),
    .b_out(b_out),
    .clk_o(clk_o),
    .led(led)
  );
  
  // system reset
  initial begin
    reset_n = 0;
    // Wait for reset
    #100;
    reset_n = 1;
  end

  // Main process for stimuli
  initial begin
    for (int file_idx = 0; file_idx < num_files; file_idx++) begin
      int stimuli_file;
      string l;
      int x, y;
      int i, r_integer, g_integer, b_integer;

      // Open the stimuli file
      stimuli_file = $fopen(stimuli_filenames[file_idx], "r");
      if (stimuli_file == 0) begin
        $display("Failed to open %s", stimuli_filenames[file_idx]);
        $finish;
      end
      $fgets(l, stimuli_file);  // read line 1 with magic number
      $fgets(l, stimuli_file);  // read line 2 with comments
      $fgets(l, stimuli_file);  // read line 3 with x, y size
      $sscanf(l, "%d %d", x_size, y_size);
      $fgets(l, stimuli_file);  // read line 4 with maximum value

      // Initialize signals
      enable_in = 3'b111;
      vs_in = 0;
      hs_in = 0;
      de_in = 0;
      r_in = 8'h00;
      g_in = 8'h00;
      b_in = 8'h00;

      // Loop for one frame
      for (y = 0; y < y_size; y++) begin
        // Set vertical sync
        if (y == 0)
          vs_in = 1;
        else
          vs_in = 0;

        // Set horizontal sync
        hs_in = 1;
        for (x = 0; x < x_blank; x++) begin
          @(negedge clk);
        end
        hs_in = 0;

        // Read one image line from file and give it to DUV
        de_in = 1;
        for (x = 0; x < x_size; x++) begin
          if ($feof(stimuli_file)) $fgets(l, stimuli_file);
          $fscanf(stimuli_file, "%d %d %d\n", r_integer, g_integer, b_integer);
          r_in = r_integer[7:0];
          g_in = g_integer[7:0];
          b_in = b_integer[7:0];
          
          @(negedge clk);
        end
        de_in = 0;
        r_in = 8'h00;
        g_in = 8'h00;
        b_in = 8'h00;
      end

      // Simulation for trailing clock cycles
      for (i = 0; i < trail; i++) begin
        @(negedge clk);
      end

      end_tb = 1; // signal to close response_file
      $fclose(stimuli_file);
      #20;

      // Stop simulation after last file
      if (file_idx == num_files - 1) begin
        $fatal("Simulation completed");
      end else begin
        end_tb = 0; // Reset the end_tb signal for the next file
      end
    end
  end

  // Second process to handle DUV output
  initial begin
    for (int file_idx = 0; file_idx < num_files; file_idx++) begin
      int response_file;
      string l_sim;
      int r_sim, g_sim, b_sim;

      wait (hs_out == 1);

      // Open file for output image
      response_file = $fopen(response_filenames[file_idx], "w");
      if (response_file == 0) begin
        $display("Failed to open %s", response_filenames[file_idx]);
        $finish;
      end
      $fwrite(response_file, "P3\n");       // magic number
      $fwrite(response_file, "# generated by SystemVerilog testbench\n");  // comment
      $fwrite(response_file, "%d %d\n", x_size, y_size);  // x, y size
      $fwrite(response_file, "255\n");  // maximum value

      while (end_tb != 1) begin
        @(negedge clk);
        if (de_out == 1) begin
          r_sim = r_out;
          g_sim = g_out;
          b_sim = b_out;
          $fwrite(response_file, "%d %d %d\n", r_sim, g_sim, b_sim);
        end
      end
      // Close respone file
      $fclose(response_file);
    end
  end

endmodule
