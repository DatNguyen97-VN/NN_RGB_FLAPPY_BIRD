package sigmoid_package;

const logic [7:0] sigmoid_lut [65536]= '{
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h02,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h03,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h07,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h08,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h09,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0A,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0B,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0D,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0E,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h0F,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h10,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h11,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h12,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h13,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h16,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h17,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h19,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1A,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1B,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1C,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1D,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1E,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h1F,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h20,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h21,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h22,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h23,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h26,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h27,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h28,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h29,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2A,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2B,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2C,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2D,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2E,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h2F,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h31,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h32,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h36,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h37,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h38,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h39,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3A,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3B,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3C,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3D,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3E,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h3F,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h40,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h41,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h42,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h43,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h44,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h45,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h46,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h47,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h48,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h49,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4A,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4B,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4C,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4D,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4E,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h4F,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h50,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h51,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h52,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h53,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h56,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h57,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h58,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h59,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5A,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5B,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5C,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5D,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5E,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h5F,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h60,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h61,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h62,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64
};

endpackage
